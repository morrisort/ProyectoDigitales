// -----------------------------------------------------------------------------
// 'pixelRadiationRegistersQ' Register Component
// Revision: 17
// -----------------------------------------------------------------------------
// Generated on 2018-04-27 at 19:11 (UTC) by airhdl version 2018.03.2
// -----------------------------------------------------------------------------
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" 
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE 
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE 
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE 
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR 
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF 
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS 
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN 
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) 
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE 
// POSSIBILITY OF SUCH DAMAGE.
// -----------------------------------------------------------------------------

`default_nettype none

module pixelRadiationRegistersQ_regs #(
    parameter AXI_ADDR_WIDTH                    = 32, // width of the AXI address bus
    parameter logic [31:0] BASEADDR = 32'h00000000 // the register file's system base address 
    ) (
    // Clock and Reset
    input  wire                                 axi_aclk,
    input  wire                                 axi_aresetn,

    // AXI Write Address Channel
    input  wire [AXI_ADDR_WIDTH-1:0]            s_axi_awaddr,
    input  wire [2:0]                           s_axi_awprot,
    input  wire                                 s_axi_awvalid,
    output wire                                 s_axi_awready,

    // AXI Write Data Channel
    input  wire [31:0]                          s_axi_wdata,
    input  wire [3:0]                           s_axi_wstrb,
    input  wire                                 s_axi_wvalid,
    output wire                                 s_axi_wready,


    // AXI Read Address Channel
    input  wire [AXI_ADDR_WIDTH-1:0]            s_axi_araddr,
    input  wire [2:0]                           s_axi_arprot,
    input  wire                                 s_axi_arvalid,
    output wire                                 s_axi_arready,

    // AXI Read Data Channel
    output wire [31:0]                          s_axi_rdata,
    output wire [1:0]                           s_axi_rresp,
    output wire                                 s_axi_rvalid,
    input  wire                                 s_axi_rready,

    // AXI Write Response Channel
    output wire [1:0]                           s_axi_bresp,
    output wire                                 s_axi_bvalid,
    input  wire                                 s_axi_bready,
    
    // User Ports          
    output wire upperresult_strobe, // Strobe logic for register 'upperResult' (pulsed when the register is read from the bus}
    input wire [31:0] upperresult_value, // Value of register 'upperResult', field 'value'
    output wire lowerresult_strobe, // Strobe logic for register 'lowerResult' (pulsed when the register is read from the bus}
    input wire [31:0] lowerresult_value, // Value of register 'lowerResult', field 'value'
    output wire dataqblue1_strobe, // Strobe logic for register 'dataQBlue1' (pulsed when the register is written from the bus}
    output wire [31:0] dataqblue1_value, // Value of register 'dataQBlue1', field 'value'
    output wire dataqblue2_strobe, // Strobe logic for register 'dataQBlue2' (pulsed when the register is written from the bus}
    output wire [31:0] dataqblue2_value, // Value of register 'dataQBlue2', field 'value'
    output wire dataqgreen1_strobe, // Strobe logic for register 'dataQGreen1' (pulsed when the register is written from the bus}
    output wire [31:0] dataqgreen1_value, // Value of register 'dataQGreen1', field 'value'
    output wire dataqgreen2_strobe, // Strobe logic for register 'dataQGreen2' (pulsed when the register is written from the bus}
    output wire [31:0] dataqgreen2_value, // Value of register 'dataQGreen2', field 'value'
    output wire dataqred1_strobe, // Strobe logic for register 'dataQRed1' (pulsed when the register is written from the bus}
    output wire [31:0] dataqred1_value, // Value of register 'dataQRed1', field 'value'
    output wire dataqred2_strobe, // Strobe logic for register 'dataQRed2' (pulsed when the register is written from the bus}
    output wire [31:0] dataqred2_value, // Value of register 'dataQRed2', field 'value'
    output wire command_strobe, // Strobe logic for register 'command' (pulsed when the register is written from the bus}
    output wire [31:0] command_value, // Value of register 'command', field 'value'
    output wire upperconstant_strobe, // Strobe logic for register 'upperConstant' (pulsed when the register is written from the bus}
    output wire [31:0] upperconstant_value, // Value of register 'upperConstant', field 'value'
    output wire lowerconstant_strobe, // Strobe logic for register 'lowerConstant' (pulsed when the register is written from the bus}
    output wire [31:0] lowerconstant_value // Value of register 'lowerConstant', field 'value'
    );

    // Constants
    localparam logic [1:0]                      AXI_OKAY        = 2'b00;
    localparam logic [1:0]                      AXI_DECERR      = 2'b11;

    // Registered signals
    logic                                       s_axi_awready_r;
    logic                                       s_axi_wready_r;
    logic [$bits(s_axi_awaddr)-1:0]             s_axi_awaddr_reg_r;
    logic                                       s_axi_bvalid_r;
    logic [$bits(s_axi_bresp)-1:0]              s_axi_bresp_r;
    logic                                       s_axi_arready_r;
    logic [$bits(s_axi_araddr)-1:0]             s_axi_araddr_reg_r;
    logic                                       s_axi_rvalid_r;
    logic [$bits(s_axi_rresp)-1:0]              s_axi_rresp_r;
    logic [$bits(s_axi_wdata)-1:0]              s_axi_wdata_reg_r;
    logic [$bits(s_axi_wstrb)-1:0]              s_axi_wstrb_reg_r;
    logic [$bits(s_axi_rdata)-1:0]              s_axi_rdata_r;
    
    // User-defined registers
    logic s_upperresult_strobe_r; // read strobe for register 'upperResult'
    logic [31:0] s_reg_upperresult_value_ro; // register 'upperResult', field 'value'
    logic s_lowerresult_strobe_r; // read strobe for register 'lowerResult'
    logic [31:0] s_reg_lowerresult_value_ro; // register 'lowerResult', field 'value'
    logic s_dataqblue1_strobe_r; // write strobe for register 'dataQBlue1'
    logic [31:0] s_reg_dataqblue1_value_rw_r; // register 'dataQBlue1', field 'value'
    logic s_dataqblue2_strobe_r; // write strobe for register 'dataQBlue2'
    logic [31:0] s_reg_dataqblue2_value_rw_r; // register 'dataQBlue2', field 'value'
    logic s_dataqgreen1_strobe_r; // write strobe for register 'dataQGreen1'
    logic [31:0] s_reg_dataqgreen1_value_rw_r; // register 'dataQGreen1', field 'value'
    logic s_dataqgreen2_strobe_r; // write strobe for register 'dataQGreen2'
    logic [31:0] s_reg_dataqgreen2_value_rw_r; // register 'dataQGreen2', field 'value'
    logic s_dataqred1_strobe_r; // write strobe for register 'dataQRed1'
    logic [31:0] s_reg_dataqred1_value_rw_r; // register 'dataQRed1', field 'value'
    logic s_dataqred2_strobe_r; // write strobe for register 'dataQRed2'
    logic [31:0] s_reg_dataqred2_value_rw_r; // register 'dataQRed2', field 'value'
    logic s_command_strobe_r; // write strobe for register 'command'
    logic [31:0] s_reg_command_value_rw_r; // register 'command', field 'value'
    logic s_upperconstant_strobe_r; // write strobe for register 'upperConstant'
    logic [31:0] s_reg_upperconstant_value_rw_r; // register 'upperConstant', field 'value'
    logic s_lowerconstant_strobe_r; // write strobe for register 'lowerConstant'
    logic [31:0] s_reg_lowerconstant_value_rw_r; // register 'lowerConstant', field 'value'

    //--------------------------------------------------------------------------
    // Inputs
    //
    assign s_reg_upperresult_value_ro = upperresult_value; // register 'upperResult', field 'value'
    assign s_reg_lowerresult_value_ro = lowerresult_value; // register 'lowerResult', field 'value'

    //--------------------------------------------------------------------------
    // Read-transaction FSM
    //    

    typedef enum {
        READ_IDLE,
        READ_REGISTER,
        READ_DONE
    } read_state_t;

    always_ff@(posedge axi_aclk or negedge axi_aresetn) begin: read_fsm
        read_state_t                                v_state_r;
        logic                                       v_addr_hit;
        if (~axi_aresetn) begin
            v_state_r          <= READ_IDLE;
            s_axi_arready_r    <= '0;
            s_axi_rvalid_r     <= '0;
            s_axi_rresp_r      <= '0;
            s_axi_araddr_reg_r <= '0;
            s_axi_rdata_r      <= '0;
            s_upperresult_strobe_r <= '0;
            s_lowerresult_strobe_r <= '0;
        end else begin
            // Default values:
            s_axi_arready_r <= 1'b0;
            s_upperresult_strobe_r <= '0;
            s_lowerresult_strobe_r <= '0;
            v_addr_hit           = 1'b0;

            case (v_state_r)

                // Wait for the start of a read transaction, which is 
                // initiated by the assertion of ARVALID
                READ_IDLE: begin
                    if (s_axi_arvalid) begin
                        s_axi_araddr_reg_r <= s_axi_araddr;     // save the read address
                        s_axi_arready_r    <= 1'b1;             // acknowledge the read-address
                        v_state_r          <= READ_REGISTER;
                    end
                end

                // Read from the actual storage element
                READ_REGISTER: begin
                    s_axi_rresp_r   <= AXI_OKAY;                // default value, may be overriden in case of decode error
                    s_axi_rvalid_r  <= 1'b1;
                    s_axi_rdata_r   <= '0;                      // default
                    
                    // register 'upperResult' at address offset 0x0
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::UPPERRESULT_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_upperresult_value_ro;
                        s_upperresult_strobe_r <= 1'b1;
                    end
                    // register 'lowerResult' at address offset 0x4
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::LOWERRESULT_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_lowerresult_value_ro;
                        s_lowerresult_strobe_r <= 1'b1;
                    end
                    // register 'dataQBlue1' at address offset 0x8
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQBLUE1_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_dataqblue1_value_rw_r;
                    end
                    // register 'dataQBlue2' at address offset 0xC
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQBLUE2_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_dataqblue2_value_rw_r;
                    end
                    // register 'dataQGreen1' at address offset 0x10
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQGREEN1_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_dataqgreen1_value_rw_r;
                    end
                    // register 'dataQGreen2' at address offset 0x14
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQGREEN2_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_dataqgreen2_value_rw_r;
                    end
                    // register 'dataQRed1' at address offset 0x18
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQRED1_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_dataqred1_value_rw_r;
                    end
                    // register 'dataQRed2' at address offset 0x1C
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQRED2_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_dataqred2_value_rw_r;
                    end
                    // register 'command' at address offset 0x20
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::COMMAND_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_command_value_rw_r;
                    end
                    // register 'upperConstant' at address offset 0x24
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::UPPERCONSTANT_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_upperconstant_value_rw_r;
                    end
                    // register 'lowerConstant' at address offset 0x28
                    if (s_axi_araddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::LOWERCONSTANT_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_axi_rdata_r[31:0] <= s_reg_lowerconstant_value_rw_r;
                    end
                    if (!v_addr_hit) begin
                        s_axi_rresp_r <= AXI_DECERR;
                        // pragma translate_off
                        $warning("ARADDR decode error");
                        // pragma translate_on
                    end
                    v_state_r <= READ_DONE;
                end
                // Write transaction completed, wait for master RREADY to proceed
                READ_DONE: begin
                    if (s_axi_rready) begin
                        s_axi_rvalid_r <= 1'b0;
                        v_state_r      <= READ_IDLE;
                    end
                end
            endcase
        end
    end: read_fsm

    //--------------------------------------------------------------------------
    // Write-transaction FSM
    //    

    typedef enum {
        WRITE_IDLE,
        WRITE_ADDR_FIRST,
        WRITE_DATA_FIRST,
        WRITE_UPDATE_REGISTER,
        WRITE_DONE
    } write_state_t;

    always_ff@(posedge axi_aclk or negedge axi_aresetn) begin: write_fsm
        write_state_t                               v_state_r;
        logic                                       v_addr_hit;
        if (~axi_aresetn) begin
            v_state_r                   <= WRITE_IDLE;
            s_axi_awready_r             <= 1'b0;
            s_axi_wready_r              <= 1'b0;
            s_axi_awaddr_reg_r          <= '0;
            s_axi_wdata_reg_r           <= '0;
            s_axi_wstrb_reg_r           <= '0;
            s_axi_bvalid_r              <= 1'b0;
            s_axi_bresp_r               <= '0;
                        
            s_dataqblue1_strobe_r <= '0;
            s_reg_dataqblue1_value_rw_r <= 32'b00000000000000000000000000000000;
            s_dataqblue2_strobe_r <= '0;
            s_reg_dataqblue2_value_rw_r <= 32'b00000000000000000000000000000000;
            s_dataqgreen1_strobe_r <= '0;
            s_reg_dataqgreen1_value_rw_r <= 32'b00000000000000000000000000000000;
            s_dataqgreen2_strobe_r <= '0;
            s_reg_dataqgreen2_value_rw_r <= 32'b00000000000000000000000000000000;
            s_dataqred1_strobe_r <= '0;
            s_reg_dataqred1_value_rw_r <= 32'b00000000000000000000000000000000;
            s_dataqred2_strobe_r <= '0;
            s_reg_dataqred2_value_rw_r <= 32'b00000000000000000000000000000000;
            s_command_strobe_r <= '0;
            s_reg_command_value_rw_r <= 32'b00000000000000000000000000000000;
            s_upperconstant_strobe_r <= '0;
            s_reg_upperconstant_value_rw_r <= 32'b00000000000000000000000000000000;
            s_lowerconstant_strobe_r <= '0;
            s_reg_lowerconstant_value_rw_r <= 32'b00000000000000000000000000000000;

        end else begin
            // Default values:
            s_axi_awready_r     <= 1'b0;
            s_axi_wready_r      <= 1'b0;
            s_dataqblue1_strobe_r <= '0;
            s_dataqblue2_strobe_r <= '0;
            s_dataqgreen1_strobe_r <= '0;
            s_dataqgreen2_strobe_r <= '0;
            s_dataqred1_strobe_r <= '0;
            s_dataqred2_strobe_r <= '0;
            s_command_strobe_r <= '0;
            s_upperconstant_strobe_r <= '0;
            s_lowerconstant_strobe_r <= '0;
            v_addr_hit          = 1'b0;
            // Self-clearing fields:
            case (v_state_r)

                // Wait for the start of a write transaction, which may be 
                // initiated by either of the following conditions:
                //   * assertion of both AWVALID and WVALID
                //   * assertion of AWVALID
                //   * assertion of WVALID
                WRITE_IDLE: begin
                    if (s_axi_awvalid && s_axi_wvalid) begin
                        s_axi_awaddr_reg_r <= s_axi_awaddr; // save the write-address 
                        s_axi_awready_r    <= 1'b1; // acknowledge the write-address
                        s_axi_wdata_reg_r  <= s_axi_wdata; // save the write-data
                        s_axi_wstrb_reg_r  <= s_axi_wstrb; // save the write-strobe
                        s_axi_wready_r     <= 1'b1; // acknowledge the write-data
                        v_state_r          <= WRITE_UPDATE_REGISTER;
                    end else if (s_axi_awvalid) begin
                        s_axi_awaddr_reg_r <= s_axi_awaddr; // save the write-address 
                        s_axi_awready_r    <= 1'b1; // acknowledge the write-address
                        v_state_r          <= WRITE_ADDR_FIRST;
                    end else if (s_axi_wvalid) begin
                        s_axi_wdata_reg_r <= s_axi_wdata; // save the write-data
                        s_axi_wstrb_reg_r <= s_axi_wstrb; // save the write-strobe
                        s_axi_wready_r    <= 1'b1; // acknowledge the write-data
                        v_state_r         <= WRITE_DATA_FIRST;
                    end
                end

                // Address-first write transaction: wait for the write-data
                WRITE_ADDR_FIRST: begin
                    if (s_axi_wvalid) begin
                        s_axi_wdata_reg_r <= s_axi_wdata; // save the write-data
                        s_axi_wstrb_reg_r <= s_axi_wstrb; // save the write-strobe
                        s_axi_wready_r    <= 1'b1; // acknowledge the write-data
                        v_state_r         <= WRITE_UPDATE_REGISTER;
                    end
                end

                // Data-first write transaction: wait for the write-address
                WRITE_DATA_FIRST: begin
                    if (s_axi_awvalid) begin
                        s_axi_awaddr_reg_r <= s_axi_awaddr; // save the write-address 
                        s_axi_awready_r    <= 1'b1; // acknowledge the write-address
                        v_state_r          <= WRITE_UPDATE_REGISTER;
                    end
                end

                // Update the actual storage element
                WRITE_UPDATE_REGISTER: begin
                    s_axi_bresp_r               <= AXI_OKAY; // default value, may be overriden in case of decode error
                    s_axi_bvalid_r              <= 1'b1;
                    


                    // register 'dataQBlue1' at address offset 0x8
                    if (s_axi_awaddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQBLUE1_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_dataqblue1_strobe_r <= 1'b1;
                        // field 'value':
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue1_value_rw_r[0] <= s_axi_wdata_reg_r[0]; // value[0]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue1_value_rw_r[1] <= s_axi_wdata_reg_r[1]; // value[1]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue1_value_rw_r[2] <= s_axi_wdata_reg_r[2]; // value[2]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue1_value_rw_r[3] <= s_axi_wdata_reg_r[3]; // value[3]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue1_value_rw_r[4] <= s_axi_wdata_reg_r[4]; // value[4]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue1_value_rw_r[5] <= s_axi_wdata_reg_r[5]; // value[5]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue1_value_rw_r[6] <= s_axi_wdata_reg_r[6]; // value[6]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue1_value_rw_r[7] <= s_axi_wdata_reg_r[7]; // value[7]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue1_value_rw_r[8] <= s_axi_wdata_reg_r[8]; // value[8]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue1_value_rw_r[9] <= s_axi_wdata_reg_r[9]; // value[9]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue1_value_rw_r[10] <= s_axi_wdata_reg_r[10]; // value[10]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue1_value_rw_r[11] <= s_axi_wdata_reg_r[11]; // value[11]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue1_value_rw_r[12] <= s_axi_wdata_reg_r[12]; // value[12]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue1_value_rw_r[13] <= s_axi_wdata_reg_r[13]; // value[13]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue1_value_rw_r[14] <= s_axi_wdata_reg_r[14]; // value[14]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue1_value_rw_r[15] <= s_axi_wdata_reg_r[15]; // value[15]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue1_value_rw_r[16] <= s_axi_wdata_reg_r[16]; // value[16]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue1_value_rw_r[17] <= s_axi_wdata_reg_r[17]; // value[17]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue1_value_rw_r[18] <= s_axi_wdata_reg_r[18]; // value[18]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue1_value_rw_r[19] <= s_axi_wdata_reg_r[19]; // value[19]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue1_value_rw_r[20] <= s_axi_wdata_reg_r[20]; // value[20]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue1_value_rw_r[21] <= s_axi_wdata_reg_r[21]; // value[21]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue1_value_rw_r[22] <= s_axi_wdata_reg_r[22]; // value[22]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue1_value_rw_r[23] <= s_axi_wdata_reg_r[23]; // value[23]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue1_value_rw_r[24] <= s_axi_wdata_reg_r[24]; // value[24]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue1_value_rw_r[25] <= s_axi_wdata_reg_r[25]; // value[25]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue1_value_rw_r[26] <= s_axi_wdata_reg_r[26]; // value[26]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue1_value_rw_r[27] <= s_axi_wdata_reg_r[27]; // value[27]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue1_value_rw_r[28] <= s_axi_wdata_reg_r[28]; // value[28]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue1_value_rw_r[29] <= s_axi_wdata_reg_r[29]; // value[29]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue1_value_rw_r[30] <= s_axi_wdata_reg_r[30]; // value[30]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue1_value_rw_r[31] <= s_axi_wdata_reg_r[31]; // value[31]
                        end
                    end

                    // register 'dataQBlue2' at address offset 0xC
                    if (s_axi_awaddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQBLUE2_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_dataqblue2_strobe_r <= 1'b1;
                        // field 'value':
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue2_value_rw_r[0] <= s_axi_wdata_reg_r[0]; // value[0]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue2_value_rw_r[1] <= s_axi_wdata_reg_r[1]; // value[1]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue2_value_rw_r[2] <= s_axi_wdata_reg_r[2]; // value[2]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue2_value_rw_r[3] <= s_axi_wdata_reg_r[3]; // value[3]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue2_value_rw_r[4] <= s_axi_wdata_reg_r[4]; // value[4]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue2_value_rw_r[5] <= s_axi_wdata_reg_r[5]; // value[5]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue2_value_rw_r[6] <= s_axi_wdata_reg_r[6]; // value[6]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqblue2_value_rw_r[7] <= s_axi_wdata_reg_r[7]; // value[7]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue2_value_rw_r[8] <= s_axi_wdata_reg_r[8]; // value[8]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue2_value_rw_r[9] <= s_axi_wdata_reg_r[9]; // value[9]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue2_value_rw_r[10] <= s_axi_wdata_reg_r[10]; // value[10]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue2_value_rw_r[11] <= s_axi_wdata_reg_r[11]; // value[11]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue2_value_rw_r[12] <= s_axi_wdata_reg_r[12]; // value[12]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue2_value_rw_r[13] <= s_axi_wdata_reg_r[13]; // value[13]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue2_value_rw_r[14] <= s_axi_wdata_reg_r[14]; // value[14]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqblue2_value_rw_r[15] <= s_axi_wdata_reg_r[15]; // value[15]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue2_value_rw_r[16] <= s_axi_wdata_reg_r[16]; // value[16]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue2_value_rw_r[17] <= s_axi_wdata_reg_r[17]; // value[17]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue2_value_rw_r[18] <= s_axi_wdata_reg_r[18]; // value[18]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue2_value_rw_r[19] <= s_axi_wdata_reg_r[19]; // value[19]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue2_value_rw_r[20] <= s_axi_wdata_reg_r[20]; // value[20]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue2_value_rw_r[21] <= s_axi_wdata_reg_r[21]; // value[21]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue2_value_rw_r[22] <= s_axi_wdata_reg_r[22]; // value[22]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqblue2_value_rw_r[23] <= s_axi_wdata_reg_r[23]; // value[23]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue2_value_rw_r[24] <= s_axi_wdata_reg_r[24]; // value[24]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue2_value_rw_r[25] <= s_axi_wdata_reg_r[25]; // value[25]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue2_value_rw_r[26] <= s_axi_wdata_reg_r[26]; // value[26]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue2_value_rw_r[27] <= s_axi_wdata_reg_r[27]; // value[27]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue2_value_rw_r[28] <= s_axi_wdata_reg_r[28]; // value[28]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue2_value_rw_r[29] <= s_axi_wdata_reg_r[29]; // value[29]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue2_value_rw_r[30] <= s_axi_wdata_reg_r[30]; // value[30]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqblue2_value_rw_r[31] <= s_axi_wdata_reg_r[31]; // value[31]
                        end
                    end

                    // register 'dataQGreen1' at address offset 0x10
                    if (s_axi_awaddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQGREEN1_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_dataqgreen1_strobe_r <= 1'b1;
                        // field 'value':
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen1_value_rw_r[0] <= s_axi_wdata_reg_r[0]; // value[0]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen1_value_rw_r[1] <= s_axi_wdata_reg_r[1]; // value[1]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen1_value_rw_r[2] <= s_axi_wdata_reg_r[2]; // value[2]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen1_value_rw_r[3] <= s_axi_wdata_reg_r[3]; // value[3]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen1_value_rw_r[4] <= s_axi_wdata_reg_r[4]; // value[4]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen1_value_rw_r[5] <= s_axi_wdata_reg_r[5]; // value[5]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen1_value_rw_r[6] <= s_axi_wdata_reg_r[6]; // value[6]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen1_value_rw_r[7] <= s_axi_wdata_reg_r[7]; // value[7]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen1_value_rw_r[8] <= s_axi_wdata_reg_r[8]; // value[8]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen1_value_rw_r[9] <= s_axi_wdata_reg_r[9]; // value[9]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen1_value_rw_r[10] <= s_axi_wdata_reg_r[10]; // value[10]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen1_value_rw_r[11] <= s_axi_wdata_reg_r[11]; // value[11]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen1_value_rw_r[12] <= s_axi_wdata_reg_r[12]; // value[12]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen1_value_rw_r[13] <= s_axi_wdata_reg_r[13]; // value[13]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen1_value_rw_r[14] <= s_axi_wdata_reg_r[14]; // value[14]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen1_value_rw_r[15] <= s_axi_wdata_reg_r[15]; // value[15]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen1_value_rw_r[16] <= s_axi_wdata_reg_r[16]; // value[16]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen1_value_rw_r[17] <= s_axi_wdata_reg_r[17]; // value[17]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen1_value_rw_r[18] <= s_axi_wdata_reg_r[18]; // value[18]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen1_value_rw_r[19] <= s_axi_wdata_reg_r[19]; // value[19]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen1_value_rw_r[20] <= s_axi_wdata_reg_r[20]; // value[20]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen1_value_rw_r[21] <= s_axi_wdata_reg_r[21]; // value[21]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen1_value_rw_r[22] <= s_axi_wdata_reg_r[22]; // value[22]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen1_value_rw_r[23] <= s_axi_wdata_reg_r[23]; // value[23]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen1_value_rw_r[24] <= s_axi_wdata_reg_r[24]; // value[24]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen1_value_rw_r[25] <= s_axi_wdata_reg_r[25]; // value[25]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen1_value_rw_r[26] <= s_axi_wdata_reg_r[26]; // value[26]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen1_value_rw_r[27] <= s_axi_wdata_reg_r[27]; // value[27]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen1_value_rw_r[28] <= s_axi_wdata_reg_r[28]; // value[28]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen1_value_rw_r[29] <= s_axi_wdata_reg_r[29]; // value[29]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen1_value_rw_r[30] <= s_axi_wdata_reg_r[30]; // value[30]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen1_value_rw_r[31] <= s_axi_wdata_reg_r[31]; // value[31]
                        end
                    end

                    // register 'dataQGreen2' at address offset 0x14
                    if (s_axi_awaddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQGREEN2_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_dataqgreen2_strobe_r <= 1'b1;
                        // field 'value':
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen2_value_rw_r[0] <= s_axi_wdata_reg_r[0]; // value[0]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen2_value_rw_r[1] <= s_axi_wdata_reg_r[1]; // value[1]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen2_value_rw_r[2] <= s_axi_wdata_reg_r[2]; // value[2]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen2_value_rw_r[3] <= s_axi_wdata_reg_r[3]; // value[3]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen2_value_rw_r[4] <= s_axi_wdata_reg_r[4]; // value[4]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen2_value_rw_r[5] <= s_axi_wdata_reg_r[5]; // value[5]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen2_value_rw_r[6] <= s_axi_wdata_reg_r[6]; // value[6]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqgreen2_value_rw_r[7] <= s_axi_wdata_reg_r[7]; // value[7]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen2_value_rw_r[8] <= s_axi_wdata_reg_r[8]; // value[8]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen2_value_rw_r[9] <= s_axi_wdata_reg_r[9]; // value[9]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen2_value_rw_r[10] <= s_axi_wdata_reg_r[10]; // value[10]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen2_value_rw_r[11] <= s_axi_wdata_reg_r[11]; // value[11]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen2_value_rw_r[12] <= s_axi_wdata_reg_r[12]; // value[12]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen2_value_rw_r[13] <= s_axi_wdata_reg_r[13]; // value[13]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen2_value_rw_r[14] <= s_axi_wdata_reg_r[14]; // value[14]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqgreen2_value_rw_r[15] <= s_axi_wdata_reg_r[15]; // value[15]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen2_value_rw_r[16] <= s_axi_wdata_reg_r[16]; // value[16]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen2_value_rw_r[17] <= s_axi_wdata_reg_r[17]; // value[17]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen2_value_rw_r[18] <= s_axi_wdata_reg_r[18]; // value[18]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen2_value_rw_r[19] <= s_axi_wdata_reg_r[19]; // value[19]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen2_value_rw_r[20] <= s_axi_wdata_reg_r[20]; // value[20]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen2_value_rw_r[21] <= s_axi_wdata_reg_r[21]; // value[21]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen2_value_rw_r[22] <= s_axi_wdata_reg_r[22]; // value[22]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqgreen2_value_rw_r[23] <= s_axi_wdata_reg_r[23]; // value[23]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen2_value_rw_r[24] <= s_axi_wdata_reg_r[24]; // value[24]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen2_value_rw_r[25] <= s_axi_wdata_reg_r[25]; // value[25]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen2_value_rw_r[26] <= s_axi_wdata_reg_r[26]; // value[26]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen2_value_rw_r[27] <= s_axi_wdata_reg_r[27]; // value[27]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen2_value_rw_r[28] <= s_axi_wdata_reg_r[28]; // value[28]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen2_value_rw_r[29] <= s_axi_wdata_reg_r[29]; // value[29]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen2_value_rw_r[30] <= s_axi_wdata_reg_r[30]; // value[30]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqgreen2_value_rw_r[31] <= s_axi_wdata_reg_r[31]; // value[31]
                        end
                    end

                    // register 'dataQRed1' at address offset 0x18
                    if (s_axi_awaddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQRED1_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_dataqred1_strobe_r <= 1'b1;
                        // field 'value':
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred1_value_rw_r[0] <= s_axi_wdata_reg_r[0]; // value[0]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred1_value_rw_r[1] <= s_axi_wdata_reg_r[1]; // value[1]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred1_value_rw_r[2] <= s_axi_wdata_reg_r[2]; // value[2]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred1_value_rw_r[3] <= s_axi_wdata_reg_r[3]; // value[3]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred1_value_rw_r[4] <= s_axi_wdata_reg_r[4]; // value[4]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred1_value_rw_r[5] <= s_axi_wdata_reg_r[5]; // value[5]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred1_value_rw_r[6] <= s_axi_wdata_reg_r[6]; // value[6]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred1_value_rw_r[7] <= s_axi_wdata_reg_r[7]; // value[7]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred1_value_rw_r[8] <= s_axi_wdata_reg_r[8]; // value[8]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred1_value_rw_r[9] <= s_axi_wdata_reg_r[9]; // value[9]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred1_value_rw_r[10] <= s_axi_wdata_reg_r[10]; // value[10]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred1_value_rw_r[11] <= s_axi_wdata_reg_r[11]; // value[11]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred1_value_rw_r[12] <= s_axi_wdata_reg_r[12]; // value[12]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred1_value_rw_r[13] <= s_axi_wdata_reg_r[13]; // value[13]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred1_value_rw_r[14] <= s_axi_wdata_reg_r[14]; // value[14]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred1_value_rw_r[15] <= s_axi_wdata_reg_r[15]; // value[15]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred1_value_rw_r[16] <= s_axi_wdata_reg_r[16]; // value[16]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred1_value_rw_r[17] <= s_axi_wdata_reg_r[17]; // value[17]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred1_value_rw_r[18] <= s_axi_wdata_reg_r[18]; // value[18]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred1_value_rw_r[19] <= s_axi_wdata_reg_r[19]; // value[19]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred1_value_rw_r[20] <= s_axi_wdata_reg_r[20]; // value[20]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred1_value_rw_r[21] <= s_axi_wdata_reg_r[21]; // value[21]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred1_value_rw_r[22] <= s_axi_wdata_reg_r[22]; // value[22]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred1_value_rw_r[23] <= s_axi_wdata_reg_r[23]; // value[23]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred1_value_rw_r[24] <= s_axi_wdata_reg_r[24]; // value[24]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred1_value_rw_r[25] <= s_axi_wdata_reg_r[25]; // value[25]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred1_value_rw_r[26] <= s_axi_wdata_reg_r[26]; // value[26]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred1_value_rw_r[27] <= s_axi_wdata_reg_r[27]; // value[27]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred1_value_rw_r[28] <= s_axi_wdata_reg_r[28]; // value[28]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred1_value_rw_r[29] <= s_axi_wdata_reg_r[29]; // value[29]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred1_value_rw_r[30] <= s_axi_wdata_reg_r[30]; // value[30]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred1_value_rw_r[31] <= s_axi_wdata_reg_r[31]; // value[31]
                        end
                    end

                    // register 'dataQRed2' at address offset 0x1C
                    if (s_axi_awaddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::DATAQRED2_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_dataqred2_strobe_r <= 1'b1;
                        // field 'value':
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred2_value_rw_r[0] <= s_axi_wdata_reg_r[0]; // value[0]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred2_value_rw_r[1] <= s_axi_wdata_reg_r[1]; // value[1]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred2_value_rw_r[2] <= s_axi_wdata_reg_r[2]; // value[2]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred2_value_rw_r[3] <= s_axi_wdata_reg_r[3]; // value[3]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred2_value_rw_r[4] <= s_axi_wdata_reg_r[4]; // value[4]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred2_value_rw_r[5] <= s_axi_wdata_reg_r[5]; // value[5]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred2_value_rw_r[6] <= s_axi_wdata_reg_r[6]; // value[6]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_dataqred2_value_rw_r[7] <= s_axi_wdata_reg_r[7]; // value[7]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred2_value_rw_r[8] <= s_axi_wdata_reg_r[8]; // value[8]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred2_value_rw_r[9] <= s_axi_wdata_reg_r[9]; // value[9]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred2_value_rw_r[10] <= s_axi_wdata_reg_r[10]; // value[10]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred2_value_rw_r[11] <= s_axi_wdata_reg_r[11]; // value[11]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred2_value_rw_r[12] <= s_axi_wdata_reg_r[12]; // value[12]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred2_value_rw_r[13] <= s_axi_wdata_reg_r[13]; // value[13]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred2_value_rw_r[14] <= s_axi_wdata_reg_r[14]; // value[14]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_dataqred2_value_rw_r[15] <= s_axi_wdata_reg_r[15]; // value[15]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred2_value_rw_r[16] <= s_axi_wdata_reg_r[16]; // value[16]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred2_value_rw_r[17] <= s_axi_wdata_reg_r[17]; // value[17]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred2_value_rw_r[18] <= s_axi_wdata_reg_r[18]; // value[18]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred2_value_rw_r[19] <= s_axi_wdata_reg_r[19]; // value[19]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred2_value_rw_r[20] <= s_axi_wdata_reg_r[20]; // value[20]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred2_value_rw_r[21] <= s_axi_wdata_reg_r[21]; // value[21]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred2_value_rw_r[22] <= s_axi_wdata_reg_r[22]; // value[22]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_dataqred2_value_rw_r[23] <= s_axi_wdata_reg_r[23]; // value[23]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred2_value_rw_r[24] <= s_axi_wdata_reg_r[24]; // value[24]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred2_value_rw_r[25] <= s_axi_wdata_reg_r[25]; // value[25]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred2_value_rw_r[26] <= s_axi_wdata_reg_r[26]; // value[26]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred2_value_rw_r[27] <= s_axi_wdata_reg_r[27]; // value[27]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred2_value_rw_r[28] <= s_axi_wdata_reg_r[28]; // value[28]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred2_value_rw_r[29] <= s_axi_wdata_reg_r[29]; // value[29]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred2_value_rw_r[30] <= s_axi_wdata_reg_r[30]; // value[30]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_dataqred2_value_rw_r[31] <= s_axi_wdata_reg_r[31]; // value[31]
                        end
                    end

                    // register 'command' at address offset 0x20
                    if (s_axi_awaddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::COMMAND_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_command_strobe_r <= 1'b1;
                        // field 'value':
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_command_value_rw_r[0] <= s_axi_wdata_reg_r[0]; // value[0]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_command_value_rw_r[1] <= s_axi_wdata_reg_r[1]; // value[1]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_command_value_rw_r[2] <= s_axi_wdata_reg_r[2]; // value[2]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_command_value_rw_r[3] <= s_axi_wdata_reg_r[3]; // value[3]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_command_value_rw_r[4] <= s_axi_wdata_reg_r[4]; // value[4]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_command_value_rw_r[5] <= s_axi_wdata_reg_r[5]; // value[5]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_command_value_rw_r[6] <= s_axi_wdata_reg_r[6]; // value[6]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_command_value_rw_r[7] <= s_axi_wdata_reg_r[7]; // value[7]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_command_value_rw_r[8] <= s_axi_wdata_reg_r[8]; // value[8]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_command_value_rw_r[9] <= s_axi_wdata_reg_r[9]; // value[9]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_command_value_rw_r[10] <= s_axi_wdata_reg_r[10]; // value[10]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_command_value_rw_r[11] <= s_axi_wdata_reg_r[11]; // value[11]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_command_value_rw_r[12] <= s_axi_wdata_reg_r[12]; // value[12]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_command_value_rw_r[13] <= s_axi_wdata_reg_r[13]; // value[13]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_command_value_rw_r[14] <= s_axi_wdata_reg_r[14]; // value[14]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_command_value_rw_r[15] <= s_axi_wdata_reg_r[15]; // value[15]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_command_value_rw_r[16] <= s_axi_wdata_reg_r[16]; // value[16]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_command_value_rw_r[17] <= s_axi_wdata_reg_r[17]; // value[17]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_command_value_rw_r[18] <= s_axi_wdata_reg_r[18]; // value[18]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_command_value_rw_r[19] <= s_axi_wdata_reg_r[19]; // value[19]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_command_value_rw_r[20] <= s_axi_wdata_reg_r[20]; // value[20]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_command_value_rw_r[21] <= s_axi_wdata_reg_r[21]; // value[21]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_command_value_rw_r[22] <= s_axi_wdata_reg_r[22]; // value[22]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_command_value_rw_r[23] <= s_axi_wdata_reg_r[23]; // value[23]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_command_value_rw_r[24] <= s_axi_wdata_reg_r[24]; // value[24]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_command_value_rw_r[25] <= s_axi_wdata_reg_r[25]; // value[25]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_command_value_rw_r[26] <= s_axi_wdata_reg_r[26]; // value[26]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_command_value_rw_r[27] <= s_axi_wdata_reg_r[27]; // value[27]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_command_value_rw_r[28] <= s_axi_wdata_reg_r[28]; // value[28]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_command_value_rw_r[29] <= s_axi_wdata_reg_r[29]; // value[29]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_command_value_rw_r[30] <= s_axi_wdata_reg_r[30]; // value[30]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_command_value_rw_r[31] <= s_axi_wdata_reg_r[31]; // value[31]
                        end
                    end

                    // register 'upperConstant' at address offset 0x24
                    if (s_axi_awaddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::UPPERCONSTANT_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_upperconstant_strobe_r <= 1'b1;
                        // field 'value':
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_upperconstant_value_rw_r[0] <= s_axi_wdata_reg_r[0]; // value[0]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_upperconstant_value_rw_r[1] <= s_axi_wdata_reg_r[1]; // value[1]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_upperconstant_value_rw_r[2] <= s_axi_wdata_reg_r[2]; // value[2]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_upperconstant_value_rw_r[3] <= s_axi_wdata_reg_r[3]; // value[3]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_upperconstant_value_rw_r[4] <= s_axi_wdata_reg_r[4]; // value[4]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_upperconstant_value_rw_r[5] <= s_axi_wdata_reg_r[5]; // value[5]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_upperconstant_value_rw_r[6] <= s_axi_wdata_reg_r[6]; // value[6]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_upperconstant_value_rw_r[7] <= s_axi_wdata_reg_r[7]; // value[7]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_upperconstant_value_rw_r[8] <= s_axi_wdata_reg_r[8]; // value[8]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_upperconstant_value_rw_r[9] <= s_axi_wdata_reg_r[9]; // value[9]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_upperconstant_value_rw_r[10] <= s_axi_wdata_reg_r[10]; // value[10]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_upperconstant_value_rw_r[11] <= s_axi_wdata_reg_r[11]; // value[11]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_upperconstant_value_rw_r[12] <= s_axi_wdata_reg_r[12]; // value[12]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_upperconstant_value_rw_r[13] <= s_axi_wdata_reg_r[13]; // value[13]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_upperconstant_value_rw_r[14] <= s_axi_wdata_reg_r[14]; // value[14]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_upperconstant_value_rw_r[15] <= s_axi_wdata_reg_r[15]; // value[15]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_upperconstant_value_rw_r[16] <= s_axi_wdata_reg_r[16]; // value[16]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_upperconstant_value_rw_r[17] <= s_axi_wdata_reg_r[17]; // value[17]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_upperconstant_value_rw_r[18] <= s_axi_wdata_reg_r[18]; // value[18]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_upperconstant_value_rw_r[19] <= s_axi_wdata_reg_r[19]; // value[19]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_upperconstant_value_rw_r[20] <= s_axi_wdata_reg_r[20]; // value[20]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_upperconstant_value_rw_r[21] <= s_axi_wdata_reg_r[21]; // value[21]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_upperconstant_value_rw_r[22] <= s_axi_wdata_reg_r[22]; // value[22]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_upperconstant_value_rw_r[23] <= s_axi_wdata_reg_r[23]; // value[23]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_upperconstant_value_rw_r[24] <= s_axi_wdata_reg_r[24]; // value[24]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_upperconstant_value_rw_r[25] <= s_axi_wdata_reg_r[25]; // value[25]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_upperconstant_value_rw_r[26] <= s_axi_wdata_reg_r[26]; // value[26]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_upperconstant_value_rw_r[27] <= s_axi_wdata_reg_r[27]; // value[27]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_upperconstant_value_rw_r[28] <= s_axi_wdata_reg_r[28]; // value[28]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_upperconstant_value_rw_r[29] <= s_axi_wdata_reg_r[29]; // value[29]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_upperconstant_value_rw_r[30] <= s_axi_wdata_reg_r[30]; // value[30]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_upperconstant_value_rw_r[31] <= s_axi_wdata_reg_r[31]; // value[31]
                        end
                    end

                    // register 'lowerConstant' at address offset 0x28
                    if (s_axi_awaddr_reg_r == BASEADDR + pixelRadiationRegistersQ_regs_pkg::LOWERCONSTANT_OFFSET) begin
                        v_addr_hit = 1'b1;
                        s_lowerconstant_strobe_r <= 1'b1;
                        // field 'value':
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_lowerconstant_value_rw_r[0] <= s_axi_wdata_reg_r[0]; // value[0]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_lowerconstant_value_rw_r[1] <= s_axi_wdata_reg_r[1]; // value[1]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_lowerconstant_value_rw_r[2] <= s_axi_wdata_reg_r[2]; // value[2]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_lowerconstant_value_rw_r[3] <= s_axi_wdata_reg_r[3]; // value[3]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_lowerconstant_value_rw_r[4] <= s_axi_wdata_reg_r[4]; // value[4]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_lowerconstant_value_rw_r[5] <= s_axi_wdata_reg_r[5]; // value[5]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_lowerconstant_value_rw_r[6] <= s_axi_wdata_reg_r[6]; // value[6]
                        end
                        if (s_axi_wstrb_reg_r[0]) begin
                            s_reg_lowerconstant_value_rw_r[7] <= s_axi_wdata_reg_r[7]; // value[7]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_lowerconstant_value_rw_r[8] <= s_axi_wdata_reg_r[8]; // value[8]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_lowerconstant_value_rw_r[9] <= s_axi_wdata_reg_r[9]; // value[9]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_lowerconstant_value_rw_r[10] <= s_axi_wdata_reg_r[10]; // value[10]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_lowerconstant_value_rw_r[11] <= s_axi_wdata_reg_r[11]; // value[11]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_lowerconstant_value_rw_r[12] <= s_axi_wdata_reg_r[12]; // value[12]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_lowerconstant_value_rw_r[13] <= s_axi_wdata_reg_r[13]; // value[13]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_lowerconstant_value_rw_r[14] <= s_axi_wdata_reg_r[14]; // value[14]
                        end
                        if (s_axi_wstrb_reg_r[1]) begin
                            s_reg_lowerconstant_value_rw_r[15] <= s_axi_wdata_reg_r[15]; // value[15]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_lowerconstant_value_rw_r[16] <= s_axi_wdata_reg_r[16]; // value[16]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_lowerconstant_value_rw_r[17] <= s_axi_wdata_reg_r[17]; // value[17]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_lowerconstant_value_rw_r[18] <= s_axi_wdata_reg_r[18]; // value[18]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_lowerconstant_value_rw_r[19] <= s_axi_wdata_reg_r[19]; // value[19]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_lowerconstant_value_rw_r[20] <= s_axi_wdata_reg_r[20]; // value[20]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_lowerconstant_value_rw_r[21] <= s_axi_wdata_reg_r[21]; // value[21]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_lowerconstant_value_rw_r[22] <= s_axi_wdata_reg_r[22]; // value[22]
                        end
                        if (s_axi_wstrb_reg_r[2]) begin
                            s_reg_lowerconstant_value_rw_r[23] <= s_axi_wdata_reg_r[23]; // value[23]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_lowerconstant_value_rw_r[24] <= s_axi_wdata_reg_r[24]; // value[24]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_lowerconstant_value_rw_r[25] <= s_axi_wdata_reg_r[25]; // value[25]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_lowerconstant_value_rw_r[26] <= s_axi_wdata_reg_r[26]; // value[26]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_lowerconstant_value_rw_r[27] <= s_axi_wdata_reg_r[27]; // value[27]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_lowerconstant_value_rw_r[28] <= s_axi_wdata_reg_r[28]; // value[28]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_lowerconstant_value_rw_r[29] <= s_axi_wdata_reg_r[29]; // value[29]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_lowerconstant_value_rw_r[30] <= s_axi_wdata_reg_r[30]; // value[30]
                        end
                        if (s_axi_wstrb_reg_r[3]) begin
                            s_reg_lowerconstant_value_rw_r[31] <= s_axi_wdata_reg_r[31]; // value[31]
                        end
                    end

                    if (!v_addr_hit) begin
                        s_axi_bresp_r   <= AXI_DECERR;
                        // pragma translate_off
                        $warning("AWADDR decode error");
                        // pragma translate_on
                    end
                    v_state_r <= WRITE_DONE;
                end

                // Write transaction completed, wait for master BREADY to proceed
                WRITE_DONE: begin
                    if (s_axi_bready) begin
                        s_axi_bvalid_r <= 1'b0;
                        v_state_r      <= WRITE_IDLE;
                    end
                end
            endcase


        end
    end: write_fsm

    //--------------------------------------------------------------------------
    // Outputs
    //
    assign s_axi_awready = s_axi_awready_r;
    assign s_axi_wready  = s_axi_wready_r;
    assign s_axi_bvalid  = s_axi_bvalid_r;
    assign s_axi_bresp   = s_axi_bresp_r;
    assign s_axi_arready = s_axi_arready_r;
    assign s_axi_rvalid  = s_axi_rvalid_r;
    assign s_axi_rresp   = s_axi_rresp_r;
    assign s_axi_rdata   = s_axi_rdata_r;
    
    assign upperresult_strobe = s_upperresult_strobe_r;
    assign lowerresult_strobe = s_lowerresult_strobe_r;
    assign dataqblue1_strobe = s_dataqblue1_strobe_r;
    assign dataqblue1_value = s_reg_dataqblue1_value_rw_r; // register 'dataQBlue1', field 'value'
    assign dataqblue2_strobe = s_dataqblue2_strobe_r;
    assign dataqblue2_value = s_reg_dataqblue2_value_rw_r; // register 'dataQBlue2', field 'value'
    assign dataqgreen1_strobe = s_dataqgreen1_strobe_r;
    assign dataqgreen1_value = s_reg_dataqgreen1_value_rw_r; // register 'dataQGreen1', field 'value'
    assign dataqgreen2_strobe = s_dataqgreen2_strobe_r;
    assign dataqgreen2_value = s_reg_dataqgreen2_value_rw_r; // register 'dataQGreen2', field 'value'
    assign dataqred1_strobe = s_dataqred1_strobe_r;
    assign dataqred1_value = s_reg_dataqred1_value_rw_r; // register 'dataQRed1', field 'value'
    assign dataqred2_strobe = s_dataqred2_strobe_r;
    assign dataqred2_value = s_reg_dataqred2_value_rw_r; // register 'dataQRed2', field 'value'
    assign command_strobe = s_command_strobe_r;
    assign command_value = s_reg_command_value_rw_r; // register 'command', field 'value'
    assign upperconstant_strobe = s_upperconstant_strobe_r;
    assign upperconstant_value = s_reg_upperconstant_value_rw_r; // register 'upperConstant', field 'value'
    assign lowerconstant_strobe = s_lowerconstant_strobe_r;
    assign lowerconstant_value = s_reg_lowerconstant_value_rw_r; // register 'lowerConstant', field 'value'

endmodule: pixelRadiationRegistersQ_regs

`resetall
